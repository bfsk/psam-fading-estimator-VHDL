LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.all;
ENTITY pilot_buffer_new IS
	PORT(
        real_in: IN integer;
		imag_in: IN integer;
		RESET: IN STD_LOGIC;
		CLK: IN STD_LOGIC;
        calculation_in_progress: in std_logic;
		serial_real_out: out integer;
        serial_imag_out: out integer
		);
END pilot_buffer_new;

ARCHITECTURE arch_pilot_buffer_new OF pilot_buffer_new IS

    type int_array is array(0 to 29) of integer;
    signal data_signals_real : int_array;
    signal data_signals_imag : int_array;
begin
	process(CLK, RESET, calculation_in_progress)
    begin
        if (RESET = '1') then
            data_signals_real(0) <= 0;
            data_signals_real(1) <= 0;
            data_signals_real(2) <= 0;
            data_signals_real(3) <= 0;
            data_signals_real(4) <= 0;
            data_signals_real(5) <= 0;
            data_signals_real(6) <= 0;
            data_signals_real(7) <= 0;
            data_signals_real(8) <= 0;
            data_signals_real(9) <= 0;
            data_signals_real(10) <= 0;
            data_signals_real(11) <= 0;
            data_signals_real(12) <= 0;
            data_signals_real(13) <= 0;
            data_signals_real(14) <= 0;
            data_signals_real(15) <= 0;
            data_signals_real(16) <= 0;
            data_signals_real(17) <= 0;
            data_signals_real(18) <= 0;
            data_signals_real(19) <= 0;
            data_signals_real(20) <= 0;
            data_signals_real(21) <= 0;
            data_signals_real(22) <= 0;
            data_signals_real(23) <= 0;
            data_signals_real(24) <= 0;
            data_signals_real(25) <= 0;
            data_signals_real(26) <= 0;
            data_signals_real(27) <= 0;
            data_signals_real(28) <= 0;
            data_signals_real(29) <= 0;

            data_signals_imag(0) <= 0;
            data_signals_imag(1) <= 0;
            data_signals_imag(2) <= 0;
            data_signals_imag(3) <= 0;
            data_signals_imag(4) <= 0;
            data_signals_imag(5) <= 0;
            data_signals_imag(6) <= 0;
            data_signals_imag(7) <= 0;
            data_signals_imag(8) <= 0;
            data_signals_imag(9) <= 0;
            data_signals_imag(10) <= 0;
            data_signals_imag(11) <= 0;
            data_signals_imag(12) <= 0;
            data_signals_imag(13) <= 0;
            data_signals_imag(14) <= 0;
            data_signals_imag(15) <= 0;
            data_signals_imag(16) <= 0;
            data_signals_imag(17) <= 0;
            data_signals_imag(18) <= 0;
            data_signals_imag(19) <= 0;
            data_signals_imag(20) <= 0;
            data_signals_imag(21) <= 0;
            data_signals_imag(22) <= 0;
            data_signals_imag(23) <= 0;
            data_signals_imag(24) <= 0;
            data_signals_imag(25) <= 0;
            data_signals_imag(26) <= 0;
            data_signals_imag(27) <= 0;
            data_signals_imag(28) <= 0;
            data_signals_imag(29) <= 0;

            serial_real_out <= 0;
            serial_imag_out <= 0;
        elsif(CLK'event and CLK = '1') then
            serial_real_out <= data_signals_real(29);
            serial_imag_out <= data_signals_imag(29);
            
            if(calculation_in_progress = '1') then
                data_signals_real(0) <= data_signals_real(29);
                data_signals_real(1) <= data_signals_real(0);
                data_signals_real(2) <= data_signals_real(1);
                data_signals_real(3) <= data_signals_real(2);
                data_signals_real(4) <= data_signals_real(3);
                data_signals_real(5) <= data_signals_real(4);
                data_signals_real(6) <= data_signals_real(5);
                data_signals_real(7) <= data_signals_real(6);
                data_signals_real(8) <= data_signals_real(7);
                data_signals_real(9) <= data_signals_real(8);
                data_signals_real(10) <= data_signals_real(9);
                data_signals_real(11) <= data_signals_real(10);
                data_signals_real(12) <= data_signals_real(11);
                data_signals_real(13) <= data_signals_real(12);
                data_signals_real(14) <= data_signals_real(13);
                data_signals_real(15) <= data_signals_real(14);
                data_signals_real(16) <= data_signals_real(15);
                data_signals_real(17) <= data_signals_real(16);
                data_signals_real(18) <= data_signals_real(17);
                data_signals_real(19) <= data_signals_real(18);
                data_signals_real(20) <= data_signals_real(19);
                data_signals_real(21) <= data_signals_real(20);
                data_signals_real(22) <= data_signals_real(21);
                data_signals_real(23) <= data_signals_real(22);
                data_signals_real(24) <= data_signals_real(23);
                data_signals_real(25) <= data_signals_real(24);
                data_signals_real(26) <= data_signals_real(25);
                data_signals_real(27) <= data_signals_real(26);
                data_signals_real(28) <= data_signals_real(27);
                data_signals_real(29) <= data_signals_real(28);

                data_signals_imag(0) <= data_signals_imag(29);
                data_signals_imag(1) <= data_signals_imag(0);
                data_signals_imag(2) <= data_signals_imag(1);
                data_signals_imag(3) <= data_signals_imag(2);
                data_signals_imag(4) <= data_signals_imag(3);
                data_signals_imag(5) <= data_signals_imag(4);
                data_signals_imag(6) <= data_signals_imag(5);
                data_signals_imag(7) <= data_signals_imag(6);
                data_signals_imag(8) <= data_signals_imag(7);
                data_signals_imag(9) <= data_signals_imag(8);
                data_signals_imag(10) <= data_signals_imag(9);
                data_signals_imag(11) <= data_signals_imag(10);
                data_signals_imag(12) <= data_signals_imag(11);
                data_signals_imag(13) <= data_signals_imag(12);
                data_signals_imag(14) <= data_signals_imag(13);
                data_signals_imag(15) <= data_signals_imag(14);
                data_signals_imag(16) <= data_signals_imag(15);
                data_signals_imag(17) <= data_signals_imag(16);
                data_signals_imag(18) <= data_signals_imag(17);
                data_signals_imag(19) <= data_signals_imag(18);
                data_signals_imag(20) <= data_signals_imag(19);
                data_signals_imag(21) <= data_signals_imag(20);
                data_signals_imag(22) <= data_signals_imag(21);
                data_signals_imag(23) <= data_signals_imag(22);
                data_signals_imag(24) <= data_signals_imag(23);
                data_signals_imag(25) <= data_signals_imag(24);
                data_signals_imag(26) <= data_signals_imag(25);
                data_signals_imag(27) <= data_signals_imag(26);
                data_signals_imag(28) <= data_signals_imag(27);
                data_signals_imag(29) <= data_signals_imag(28);
            else
                data_signals_real(0) <= real_in;
                data_signals_real(1) <= data_signals_real(0);
                data_signals_real(2) <= data_signals_real(1);
                data_signals_real(3) <= data_signals_real(2);
                data_signals_real(4) <= data_signals_real(3);
                data_signals_real(5) <= data_signals_real(4);
                data_signals_real(6) <= data_signals_real(5);
                data_signals_real(7) <= data_signals_real(6);
                data_signals_real(8) <= data_signals_real(7);
                data_signals_real(9) <= data_signals_real(8);
                data_signals_real(10) <= data_signals_real(9);
                data_signals_real(11) <= data_signals_real(10);
                data_signals_real(12) <= data_signals_real(11);
                data_signals_real(13) <= data_signals_real(12);
                data_signals_real(14) <= data_signals_real(13);
                data_signals_real(15) <= data_signals_real(14);
                data_signals_real(16) <= data_signals_real(15);
                data_signals_real(17) <= data_signals_real(16);
                data_signals_real(18) <= data_signals_real(17);
                data_signals_real(19) <= data_signals_real(18);
                data_signals_real(20) <= data_signals_real(19);
                data_signals_real(21) <= data_signals_real(20);
                data_signals_real(22) <= data_signals_real(21);
                data_signals_real(23) <= data_signals_real(22);
                data_signals_real(24) <= data_signals_real(23);
                data_signals_real(25) <= data_signals_real(24);
                data_signals_real(26) <= data_signals_real(25);
                data_signals_real(27) <= data_signals_real(26);
                data_signals_real(28) <= data_signals_real(27);
                data_signals_real(29) <= data_signals_real(28);

                data_signals_imag(0) <= imag_in;
                data_signals_imag(1) <= data_signals_imag(0);
                data_signals_imag(2) <= data_signals_imag(1);
                data_signals_imag(3) <= data_signals_imag(2);
                data_signals_imag(4) <= data_signals_imag(3);
                data_signals_imag(5) <= data_signals_imag(4);
                data_signals_imag(6) <= data_signals_imag(5);
                data_signals_imag(7) <= data_signals_imag(6);
                data_signals_imag(8) <= data_signals_imag(7);
                data_signals_imag(9) <= data_signals_imag(8);
                data_signals_imag(10) <= data_signals_imag(9);
                data_signals_imag(11) <= data_signals_imag(10);
                data_signals_imag(12) <= data_signals_imag(11);
                data_signals_imag(13) <= data_signals_imag(12);
                data_signals_imag(14) <= data_signals_imag(13);
                data_signals_imag(15) <= data_signals_imag(14);
                data_signals_imag(16) <= data_signals_imag(15);
                data_signals_imag(17) <= data_signals_imag(16);
                data_signals_imag(18) <= data_signals_imag(17);
                data_signals_imag(19) <= data_signals_imag(18);
                data_signals_imag(20) <= data_signals_imag(19);
                data_signals_imag(21) <= data_signals_imag(20);
                data_signals_imag(22) <= data_signals_imag(21);
                data_signals_imag(23) <= data_signals_imag(22);
                data_signals_imag(24) <= data_signals_imag(23);
                data_signals_imag(25) <= data_signals_imag(24);
                data_signals_imag(26) <= data_signals_imag(25);
                data_signals_imag(27) <= data_signals_imag(26);
                data_signals_imag(28) <= data_signals_imag(27);
                data_signals_imag(29) <= data_signals_imag(28);
            end if;
        end if;

    end process;

END ARCHITECTURE;