LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.all;

ENTITY sinc_coefficients IS
	PORT(
		index_of_symbol: IN std_logic_vector(3 downto 0);		  
		sinc_m14 : OUT integer;
	  	sinc_m13 : OUT integer;
	  	sinc_m12 : OUT integer;
	  	sinc_m11 : OUT integer;
	  	sinc_m10 : OUT integer;
	  	sinc_m9 : OUT integer;
	  	sinc_m8 : OUT integer;
	  	sinc_m7 : OUT integer;
	  	sinc_m6 : OUT integer;
	  	sinc_m5 : OUT integer;
	  	sinc_m4 : OUT integer;
	 	sinc_m3 : OUT integer;
	 	sinc_m2 : OUT integer;
		sinc_m1 : OUT integer;
		sinc_0 : OUT integer;
		sinc_1 : OUT integer;
		sinc_2 : OUT integer;
		sinc_3 : OUT integer;
		sinc_4 : OUT integer;
	  	sinc_5 : OUT integer;
	  	sinc_6 : OUT integer;
	 	sinc_7 : OUT integer;
	 	sinc_8 : OUT integer;
	 	sinc_9 : OUT integer;
		sinc_10 : OUT integer;
	 	sinc_11 : OUT integer;
	 	sinc_12 : OUT integer;
	 	sinc_13 : OUT integer;
	 	sinc_14 : OUT integer;
	 	sinc_15 : OUT integer
		);
END sinc_coefficients;

ARCHITECTURE arch_sinc_coefficients OF sinc_coefficients IS
begin

process(index_of_symbol) is
begin
	case index_of_symbol is
                when "0010"=>
        sinc_m14 <= 4704;
        sinc_m13 <= -5064;
        sinc_m12 <= 5484;
        sinc_m11 <= -5980;
        sinc_m10 <= 6574;
        sinc_m9 <= -7299;
        sinc_m8 <= 8204;
        sinc_m7 <= -9365;
        sinc_m6 <= 10908;
        sinc_m5 <= -13061;
        sinc_m4 <= 16273;
        sinc_m3 <= -21580;
        sinc_m2 <= 32022;
        sinc_m1 <= -62044;
        sinc_0 <= 992705;
        sinc_1 <= 70907;
        sinc_2 <= -34231;
        sinc_3 <= 22561;
        sinc_4 <= -16825;
        sinc_5 <= 13414;
        sinc_6 <= -11153;
        sinc_7 <= 9545;
        sinc_8 <= -8342;
        sinc_9 <= 7408;
        sinc_10 <= -6662;
        sinc_11 <= 6053;
        sinc_12 <= -5545;
        sinc_13 <= 5117;
        sinc_14 <= -4749;
        sinc_15 <= 4431;

when "0011"=>
        sinc_m14 <= 9160;
        sinc_m13 <= -9857;
        sinc_m12 <= 10670;
        sinc_m11 <= -11628;
        sinc_m10 <= 12776;
        sinc_m9 <= -14175;
        sinc_m8 <= 15918;
        sinc_m7 <= -18149;
        sinc_m6 <= 21108;
        sinc_m5 <= -25221;
        sinc_m4 <= 31322;
        sinc_m3 <= -41319;
        sinc_m2 <= 60688;
        sinc_m1 <= -114236;
        sinc_0 <= 971012;
        sinc_1 <= 149386;
        sinc_2 <= -69358;
        sinc_3 <= 45163;
        sinc_4 <= -33483;
        sinc_5 <= 26603;
        sinc_6 <= -22068;
        sinc_7 <= 18854;
        sinc_8 <= -16457;
        sinc_9 <= 14601;
        sinc_10 <= -13121;
        sinc_11 <= 11914;
        sinc_12 <= -10910;
        sinc_13 <= 10062;
        sinc_14 <= -9336;
        sinc_15 <= 8708;

when "0100"=>
        sinc_m14 <= 13175;
        sinc_m13 <= -14174;
        sinc_m12 <= 15335;
        sinc_m11 <= -16705;
        sinc_m10 <= 18342;
        sinc_m9 <= -20336;
        sinc_m8 <= 22816;
        sinc_m7 <= -25985;
        sinc_m6 <= 30177;
        sinc_m5 <= -35980;
        sinc_m4 <= 44547;
        sinc_m3 <= -58468;
        sinc_m2 <= 85044;
        sinc_m1 <= -155914;
        sinc_0 <= 935489;
        sinc_1 <= 233872;
        sinc_2 <= -103943;
        sinc_3 <= 66820;
        sinc_4 <= -49236;
        sinc_5 <= 38978;
        sinc_6 <= -32258;
        sinc_7 <= 27514;
        sinc_8 <= -23986;
        sinc_9 <= 21261;
        sinc_10 <= -19091;
        sinc_11 <= 17323;
        sinc_12 <= -15855;
        sinc_13 <= 14617;
        sinc_14 <= -13557;
        sinc_15 <= 12641;

when "0101"=>
        sinc_m14 <= 16580;
        sinc_m13 <= -17830;
        sinc_m12 <= 19283;
        sinc_m11 <= -20995;
        sinc_m10 <= 23040;
        sinc_m9 <= -25527;
        sinc_m8 <= 28614;
        sinc_m7 <= -32552;
        sinc_m6 <= 37747;
        sinc_m5 <= -44914;
        sinc_m4 <= 55441;
        sinc_m3 <= -72413;
        sinc_m2 <= 104360;
        sinc_m1 <= -186750;
        sinc_0 <= 887063;
        sinc_1 <= 322568;
        sinc_2 <= -136471;
        sinc_3 <= 86542;
        sinc_4 <= -63361;
        sinc_5 <= 49975;
        sinc_6 <= -41258;
        sinc_7 <= 35131;
        sinc_8 <= -30588;
        sinc_9 <= 27085;
        sinc_10 <= -24303;
        sinc_11 <= 22038;
        sinc_12 <= -20160;
        sinc_13 <= 18577;
        sinc_14 <= -17224;
        sinc_15 <= 16055;

when "0110"=>
        sinc_m14 <= 19232;
        sinc_m13 <= -20674;
        sinc_m12 <= 22351;
        sinc_m11 <= -24323;
        sinc_m10 <= 26677;
        sinc_m9 <= -29535;
        sinc_m8 <= 33079;
        sinc_m7 <= -37590;
        sinc_m6 <= 43525;
        sinc_m5 <= -51687;
        sinc_m4 <= 63614;
        sinc_m3 <= -82699;
        sinc_m2 <= 118141;
        sinc_m1 <= -206748;
        sinc_0 <= 826993;
        sinc_1 <= 413496;
        sinc_2 <= -165398;
        sinc_3 <= 103374;
        sinc_4 <= -75181;
        sinc_5 <= 59070;
        sinc_6 <= -48646;
        sinc_7 <= 41349;
        sinc_8 <= -35956;
        sinc_9 <= 31807;
        sinc_10 <= -28517;
        sinc_11 <= 25843;
        sinc_12 <= -23628;
        sinc_13 <= 21762;
        sinc_14 <= -20170;
        sinc_15 <= 18795;

when "0111"=>
        sinc_m14 <= 21022;
        sinc_m13 <= -22591;
        sinc_m12 <= 24413;
        sinc_m11 <= -26555;
        sinc_m10 <= 29108;
        sinc_m9 <= -32205;
        sinc_m8 <= 36039;
        sinc_m7 <= -40909;
        sinc_m6 <= 47301;
        sinc_m5 <= -56061;
        sinc_m4 <= 68802;
        sinc_m3 <= -89038;
        sinc_m2 <= 126137;
        sinc_m1 <= -216236;
        sinc_0 <= 756826;
        sinc_1 <= 504551;
        sinc_2 <= -189206;
        sinc_3 <= 116434;
        sinc_4 <= -84091;
        sinc_5 <= 65811;
        sinc_6 <= -54059;
        sinc_7 <= 45868;
        sinc_8 <= -39832;
        sinc_9 <= 35201;
        sinc_10 <= -31534;
        sinc_11 <= 28559;
        sinc_12 <= -26097;
        sinc_13 <= 24026;
        sinc_14 <= -22259;
        sinc_15 <= 20734;

when "1000"=>
        sinc_m14 <= 21882;
        sinc_m13 <= -23507;
        sinc_m12 <= 25393;
        sinc_m11 <= -27607;
        sinc_m10 <= 30245;
        sinc_m9 <= -33440;
        sinc_m8 <= 37389;
        sinc_m7 <= -42397;
        sinc_m6 <= 48953;
        sinc_m5 <= -57908;
        sinc_m4 <= 70873;
        sinc_m3 <= -91317;
        sinc_m2 <= 128337;
        sinc_m1 <= -215840;
        sinc_0 <= 678356;
        sinc_1 <= 593561;
        sinc_2 <= -206456;
        sinc_3 <= 124960;
        sinc_4 <= -89594;
        sinc_5 <= 69830;
        sinc_6 <= -57210;
        sinc_7 <= 48454;
        sinc_8 <= -42022;
        sinc_9 <= 37097;
        sinc_10 <= -33206;
        sinc_11 <= 30053;
        sinc_12 <= -27447;
        sinc_13 <= 25257;
        sinc_14 <= -23391;
        sinc_15 <= 21782;

when "1001"=>
        sinc_m14 <= 21782;
        sinc_m13 <= -23391;
        sinc_m12 <= 25257;
        sinc_m11 <= -27447;
        sinc_m10 <= 30053;
        sinc_m9 <= -33206;
        sinc_m8 <= 37097;
        sinc_m7 <= -42022;
        sinc_m6 <= 48454;
        sinc_m5 <= -57210;
        sinc_m4 <= 69830;
        sinc_m3 <= -89594;
        sinc_m2 <= 124960;
        sinc_m1 <= -206456;
        sinc_0 <= 593561;
        sinc_1 <= 678356;
        sinc_2 <= -215840;
        sinc_3 <= 128337;
        sinc_4 <= -91317;
        sinc_5 <= 70873;
        sinc_6 <= -57908;
        sinc_7 <= 48953;
        sinc_8 <= -42397;
        sinc_9 <= 37389;
        sinc_10 <= -33440;
        sinc_11 <= 30245;
        sinc_12 <= -27607;
        sinc_13 <= 25393;
        sinc_14 <= -23507;
        sinc_15 <= 21882;

when "1010"=>
        sinc_m14 <= 20734;
        sinc_m13 <= -22259;
        sinc_m12 <= 24026;
        sinc_m11 <= -26097;
        sinc_m10 <= 28559;
        sinc_m9 <= -31534;
        sinc_m8 <= 35201;
        sinc_m7 <= -39832;
        sinc_m6 <= 45868;
        sinc_m5 <= -54059;
        sinc_m4 <= 65811;
        sinc_m3 <= -84091;
        sinc_m2 <= 116434;
        sinc_m1 <= -189206;
        sinc_0 <= 504551;
        sinc_1 <= 756826;
        sinc_2 <= -216236;
        sinc_3 <= 126137;
        sinc_4 <= -89038;
        sinc_5 <= 68802;
        sinc_6 <= -56061;
        sinc_7 <= 47301;
        sinc_8 <= -40909;
        sinc_9 <= 36039;
        sinc_10 <= -32205;
        sinc_11 <= 29108;
        sinc_12 <= -26555;
        sinc_13 <= 24413;
        sinc_14 <= -22591;
        sinc_15 <= 21022;

when "1011"=>
        sinc_m14 <= 18795;
        sinc_m13 <= -20170;
        sinc_m12 <= 21762;
        sinc_m11 <= -23628;
        sinc_m10 <= 25843;
        sinc_m9 <= -28517;
        sinc_m8 <= 31807;
        sinc_m7 <= -35956;
        sinc_m6 <= 41349;
        sinc_m5 <= -48646;
        sinc_m4 <= 59070;
        sinc_m3 <= -75181;
        sinc_m2 <= 103374;
        sinc_m1 <= -165398;
        sinc_0 <= 413496;
        sinc_1 <= 826993;
        sinc_2 <= -206748;
        sinc_3 <= 118141;
        sinc_4 <= -82699;
        sinc_5 <= 63614;
        sinc_6 <= -51687;
        sinc_7 <= 43525;
        sinc_8 <= -37590;
        sinc_9 <= 33079;
        sinc_10 <= -29535;
        sinc_11 <= 26677;
        sinc_12 <= -24323;
        sinc_13 <= 22351;
        sinc_14 <= -20674;
        sinc_15 <= 19232;

when "1100"=>
        sinc_m14 <= 16055;
        sinc_m13 <= -17224;
        sinc_m12 <= 18577;
        sinc_m11 <= -20160;
        sinc_m10 <= 22038;
        sinc_m9 <= -24303;
        sinc_m8 <= 27085;
        sinc_m7 <= -30588;
        sinc_m6 <= 35131;
        sinc_m5 <= -41258;
        sinc_m4 <= 49975;
        sinc_m3 <= -63361;
        sinc_m2 <= 86542;
        sinc_m1 <= -136471;
        sinc_0 <= 322568;
        sinc_1 <= 887063;
        sinc_2 <= -186750;
        sinc_3 <= 104360;
        sinc_4 <= -72413;
        sinc_5 <= 55441;
        sinc_6 <= -44914;
        sinc_7 <= 37747;
        sinc_8 <= -32552;
        sinc_9 <= 28614;
        sinc_10 <= -25527;
        sinc_11 <= 23040;
        sinc_12 <= -20995;
        sinc_13 <= 19283;
        sinc_14 <= -17830;
        sinc_15 <= 16580;

when "1101"=>
        sinc_m14 <= 12641;
        sinc_m13 <= -13557;
        sinc_m12 <= 14617;
        sinc_m11 <= -15855;
        sinc_m10 <= 17323;
        sinc_m9 <= -19091;
        sinc_m8 <= 21261;
        sinc_m7 <= -23986;
        sinc_m6 <= 27514;
        sinc_m5 <= -32258;
        sinc_m4 <= 38978;
        sinc_m3 <= -49236;
        sinc_m2 <= 66820;
        sinc_m1 <= -103943;
        sinc_0 <= 233872;
        sinc_1 <= 935489;
        sinc_2 <= -155914;
        sinc_3 <= 85044;
        sinc_4 <= -58468;
        sinc_5 <= 44547;
        sinc_6 <= -35980;
        sinc_7 <= 30177;
        sinc_8 <= -25985;
        sinc_9 <= 22816;
        sinc_10 <= -20336;
        sinc_11 <= 18342;
        sinc_12 <= -16705;
        sinc_13 <= 15335;
        sinc_14 <= -14174;
        sinc_15 <= 13175;

when "1110"=>
        sinc_m14 <= 8708;
        sinc_m13 <= -9336;
        sinc_m12 <= 10062;
        sinc_m11 <= -10910;
        sinc_m10 <= 11914;
        sinc_m9 <= -13121;
        sinc_m8 <= 14601;
        sinc_m7 <= -16457;
        sinc_m6 <= 18854;
        sinc_m5 <= -22068;
        sinc_m4 <= 26603;
        sinc_m3 <= -33483;
        sinc_m2 <= 45163;
        sinc_m1 <= -69358;
        sinc_0 <= 149386;
        sinc_1 <= 971012;
        sinc_2 <= -114236;
        sinc_3 <= 60688;
        sinc_4 <= -41319;
        sinc_5 <= 31322;
        sinc_6 <= -25221;
        sinc_7 <= 21108;
        sinc_8 <= -18149;
        sinc_9 <= 15918;
        sinc_10 <= -14175;
        sinc_11 <= 12776;
        sinc_12 <= -11628;
        sinc_13 <= 10670;
        sinc_14 <= -9857;
        sinc_15 <= 9160;

when "1111"=>
        sinc_m14 <= 4431;
        sinc_m13 <= -4749;
        sinc_m12 <= 5117;
        sinc_m11 <= -5545;
        sinc_m10 <= 6053;
        sinc_m9 <= -6662;
        sinc_m8 <= 7408;
        sinc_m7 <= -8342;
        sinc_m6 <= 9545;
        sinc_m5 <= -11153;
        sinc_m4 <= 13414;
        sinc_m3 <= -16825;
        sinc_m2 <= 22561;
        sinc_m1 <= -34231;
        sinc_0 <= 70907;
        sinc_1 <= 992705;
        sinc_2 <= -62044;
        sinc_3 <= 32022;
        sinc_4 <= -21580;
        sinc_5 <= 16273;
        sinc_6 <= -13061;
        sinc_7 <= 10908;
        sinc_8 <= -9365;
        sinc_9 <= 8204;
        sinc_10 <= -7299;
        sinc_11 <= 6574;
        sinc_12 <= -5980;
        sinc_13 <= 5484;
        sinc_14 <= -5064;
        sinc_15 <= 4704;
  when others=> -- 0 and others
			  sinc_m14 <= 0;
			  sinc_m13 <= 0;
			  sinc_m12 <= 0;
			  sinc_m11 <= 0;
			  sinc_m10 <= 0;
			  sinc_m9 <= 0;
			  sinc_m8 <= 0;
			  sinc_m7 <= 0;
			  sinc_m6 <= 0;
			  sinc_m5 <= 0;
			  sinc_m4 <= 0;
			  sinc_m3 <= 0;
			  sinc_m2 <= 0;
			  sinc_m1 <= 0;
			  sinc_0 <= 0;
			  sinc_1 <= 0;
			  sinc_2 <= 0;
			  sinc_3 <= 0;
			  sinc_4 <= 0;
			  sinc_5 <= 0;
			  sinc_6 <= 0;
			  sinc_7 <= 0;
			  sinc_8 <= 0;
			  sinc_9 <= 0;
			  sinc_10 <= 0;
			  sinc_11 <= 0;
			  sinc_12 <= 0;
			  sinc_13 <= 0;
			  sinc_14 <= 0;
			  sinc_15 <= 0;


	end case;
end process;
END ARCHITECTURE;